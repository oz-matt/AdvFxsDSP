//-----------------------------------------------------------------------------
// Automatically generated Verilog code for non-primitive component
// Design1_1.v
//-----------------------------------------------------------------------------
`timescale 1ns/10ps
//-----------------------------------------------------------------------------
// declare Design1_1 module
//-----------------------------------------------------------------------------
module Design1_1
(
    input ce1,
    input clk,
    input [31 : 0] dp1,
    output [31 : 0] dp2,
    input rst
);


//-------------------------------------------------------------------------
// declare signals
//-------------------------------------------------------------------------
wire [31 : 0] F1_dataOut;
//-------------------------------------------------------------------------
